`include "utils.svh"

module system_tb();

    test_program test();
    test_harness `TH();

endmodule
